interface wdtif;
logic wdt_intr;
endinterface
