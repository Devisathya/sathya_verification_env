library verilog;
use verilog.vl_types.all;
entity top1_sv_unit is
end top1_sv_unit;
