library verilog;
use verilog.vl_types.all;
entity wdtif is
end wdtif;
